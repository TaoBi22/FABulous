//NumberOfConfigBits:280
module RAM_IO_switch_matrix (N1END0, N1END1, N1END2, N1END3, N2MID0, N2MID1, N2MID2, N2MID3, N2MID4, N2MID5, N2MID6, N2MID7, N2END0, N2END1, N2END2, N2END3, N2END4, N2END5, N2END6, N2END7, N4END0, N4END1, N4END2, N4END3, E1END0, E1END1, E1END2, E1END3, E2MID0, E2MID1, E2MID2, E2MID3, E2MID4, E2MID5, E2MID6, E2MID7, E2END0, E2END1, E2END2, E2END3, E2END4, E2END5, E2END6, E2END7, EE4END0, EE4END1, EE4END2, EE4END3, EE4END4, EE4END5, EE4END6, EE4END7, EE4END8, EE4END9, EE4END10, EE4END11, EE4END12, EE4END13, EE4END14, EE4END15, E6END0, E6END1, E6END2, E6END3, E6END4, E6END5, E6END6, E6END7, E6END8, E6END9, E6END10, E6END11, S1END0, S1END1, S1END2, S1END3, S2MID0, S2MID1, S2MID2, S2MID3, S2MID4, S2MID5, S2MID6, S2MID7, S2END0, S2END1, S2END2, S2END3, S2END4, S2END5, S2END6, S2END7, S4END0, S4END1, S4END2, S4END3, RAM2FAB_D0_O0, RAM2FAB_D0_O1, RAM2FAB_D0_O2, RAM2FAB_D0_O3, RAM2FAB_D1_O0, RAM2FAB_D1_O1, RAM2FAB_D1_O2, RAM2FAB_D1_O3, RAM2FAB_D2_O0, RAM2FAB_D2_O1, RAM2FAB_D2_O2, RAM2FAB_D2_O3, RAM2FAB_D3_O0, RAM2FAB_D3_O1, RAM2FAB_D3_O2, RAM2FAB_D3_O3, J_NS4_END0, J_NS4_END1, J_NS4_END2, J_NS4_END3, J_NS4_END4, J_NS4_END5, J_NS4_END6, J_NS4_END7, J_NS4_END8, J_NS4_END9, J_NS4_END10, J_NS4_END11, J_NS4_END12, J_NS4_END13, J_NS4_END14, J_NS4_END15, J_NS2_END0, J_NS2_END1, J_NS2_END2, J_NS2_END3, J_NS2_END4, J_NS2_END5, J_NS2_END6, J_NS2_END7, J_NS1_END0, J_NS1_END1, J_NS1_END2, J_NS1_END3, N1BEG0, N1BEG1, N1BEG2, N1BEG3, N2BEG0, N2BEG1, N2BEG2, N2BEG3, N2BEG4, N2BEG5, N2BEG6, N2BEG7, N2BEGb0, N2BEGb1, N2BEGb2, N2BEGb3, N2BEGb4, N2BEGb5, N2BEGb6, N2BEGb7, N4BEG0, N4BEG1, N4BEG2, N4BEG3, S1BEG0, S1BEG1, S1BEG2, S1BEG3, S2BEG0, S2BEG1, S2BEG2, S2BEG3, S2BEG4, S2BEG5, S2BEG6, S2BEG7, S2BEGb0, S2BEGb1, S2BEGb2, S2BEGb3, S2BEGb4, S2BEGb5, S2BEGb6, S2BEGb7, S4BEG0, S4BEG1, S4BEG2, S4BEG3, W1BEG0, W1BEG1, W1BEG2, W1BEG3, W2BEG0, W2BEG1, W2BEG2, W2BEG3, W2BEG4, W2BEG5, W2BEG6, W2BEG7, W2BEGb0, W2BEGb1, W2BEGb2, W2BEGb3, W2BEGb4, W2BEGb5, W2BEGb6, W2BEGb7, WW4BEG0, WW4BEG1, WW4BEG2, WW4BEG3, WW4BEG4, WW4BEG5, WW4BEG6, WW4BEG7, WW4BEG8, WW4BEG9, WW4BEG10, WW4BEG11, WW4BEG12, WW4BEG13, WW4BEG14, WW4BEG15, W6BEG0, W6BEG1, W6BEG2, W6BEG3, W6BEG4, W6BEG5, W6BEG6, W6BEG7, W6BEG8, W6BEG9, W6BEG10, W6BEG11, FAB2RAM_D0_I0, FAB2RAM_D0_I1, FAB2RAM_D0_I2, FAB2RAM_D0_I3, FAB2RAM_D1_I0, FAB2RAM_D1_I1, FAB2RAM_D1_I2, FAB2RAM_D1_I3, FAB2RAM_D2_I0, FAB2RAM_D2_I1, FAB2RAM_D2_I2, FAB2RAM_D2_I3, FAB2RAM_D3_I0, FAB2RAM_D3_I1, FAB2RAM_D3_I2, FAB2RAM_D3_I3, FAB2RAM_A0_I0, FAB2RAM_A0_I1, FAB2RAM_A0_I2, FAB2RAM_A0_I3, FAB2RAM_A1_I0, FAB2RAM_A1_I1, FAB2RAM_A1_I2, FAB2RAM_A1_I3, FAB2RAM_C_I0, FAB2RAM_C_I1, FAB2RAM_C_I2, FAB2RAM_C_I3, J_NS4_BEG0, J_NS4_BEG1, J_NS4_BEG2, J_NS4_BEG3, J_NS4_BEG4, J_NS4_BEG5, J_NS4_BEG6, J_NS4_BEG7, J_NS4_BEG8, J_NS4_BEG9, J_NS4_BEG10, J_NS4_BEG11, J_NS4_BEG12, J_NS4_BEG13, J_NS4_BEG14, J_NS4_BEG15, J_NS2_BEG0, J_NS2_BEG1, J_NS2_BEG2, J_NS2_BEG3, J_NS2_BEG4, J_NS2_BEG5, J_NS2_BEG6, J_NS2_BEG7, J_NS1_BEG0, J_NS1_BEG1, J_NS1_BEG2, J_NS1_BEG3, ConfigBits, ConfigBits_N);
	parameter NoConfigBits = 280;
	 // switch matrix inputs
	input N1END0;
	input N1END1;
	input N1END2;
	input N1END3;
	input N2MID0;
	input N2MID1;
	input N2MID2;
	input N2MID3;
	input N2MID4;
	input N2MID5;
	input N2MID6;
	input N2MID7;
	input N2END0;
	input N2END1;
	input N2END2;
	input N2END3;
	input N2END4;
	input N2END5;
	input N2END6;
	input N2END7;
	input N4END0;
	input N4END1;
	input N4END2;
	input N4END3;
	input E1END0;
	input E1END1;
	input E1END2;
	input E1END3;
	input E2MID0;
	input E2MID1;
	input E2MID2;
	input E2MID3;
	input E2MID4;
	input E2MID5;
	input E2MID6;
	input E2MID7;
	input E2END0;
	input E2END1;
	input E2END2;
	input E2END3;
	input E2END4;
	input E2END5;
	input E2END6;
	input E2END7;
	input EE4END0;
	input EE4END1;
	input EE4END2;
	input EE4END3;
	input EE4END4;
	input EE4END5;
	input EE4END6;
	input EE4END7;
	input EE4END8;
	input EE4END9;
	input EE4END10;
	input EE4END11;
	input EE4END12;
	input EE4END13;
	input EE4END14;
	input EE4END15;
	input E6END0;
	input E6END1;
	input E6END2;
	input E6END3;
	input E6END4;
	input E6END5;
	input E6END6;
	input E6END7;
	input E6END8;
	input E6END9;
	input E6END10;
	input E6END11;
	input S1END0;
	input S1END1;
	input S1END2;
	input S1END3;
	input S2MID0;
	input S2MID1;
	input S2MID2;
	input S2MID3;
	input S2MID4;
	input S2MID5;
	input S2MID6;
	input S2MID7;
	input S2END0;
	input S2END1;
	input S2END2;
	input S2END3;
	input S2END4;
	input S2END5;
	input S2END6;
	input S2END7;
	input S4END0;
	input S4END1;
	input S4END2;
	input S4END3;
	input RAM2FAB_D0_O0;
	input RAM2FAB_D0_O1;
	input RAM2FAB_D0_O2;
	input RAM2FAB_D0_O3;
	input RAM2FAB_D1_O0;
	input RAM2FAB_D1_O1;
	input RAM2FAB_D1_O2;
	input RAM2FAB_D1_O3;
	input RAM2FAB_D2_O0;
	input RAM2FAB_D2_O1;
	input RAM2FAB_D2_O2;
	input RAM2FAB_D2_O3;
	input RAM2FAB_D3_O0;
	input RAM2FAB_D3_O1;
	input RAM2FAB_D3_O2;
	input RAM2FAB_D3_O3;
	input J_NS4_END0;
	input J_NS4_END1;
	input J_NS4_END2;
	input J_NS4_END3;
	input J_NS4_END4;
	input J_NS4_END5;
	input J_NS4_END6;
	input J_NS4_END7;
	input J_NS4_END8;
	input J_NS4_END9;
	input J_NS4_END10;
	input J_NS4_END11;
	input J_NS4_END12;
	input J_NS4_END13;
	input J_NS4_END14;
	input J_NS4_END15;
	input J_NS2_END0;
	input J_NS2_END1;
	input J_NS2_END2;
	input J_NS2_END3;
	input J_NS2_END4;
	input J_NS2_END5;
	input J_NS2_END6;
	input J_NS2_END7;
	input J_NS1_END0;
	input J_NS1_END1;
	input J_NS1_END2;
	input J_NS1_END3;
	output N1BEG0;
	output N1BEG1;
	output N1BEG2;
	output N1BEG3;
	output N2BEG0;
	output N2BEG1;
	output N2BEG2;
	output N2BEG3;
	output N2BEG4;
	output N2BEG5;
	output N2BEG6;
	output N2BEG7;
	output N2BEGb0;
	output N2BEGb1;
	output N2BEGb2;
	output N2BEGb3;
	output N2BEGb4;
	output N2BEGb5;
	output N2BEGb6;
	output N2BEGb7;
	output N4BEG0;
	output N4BEG1;
	output N4BEG2;
	output N4BEG3;
	output S1BEG0;
	output S1BEG1;
	output S1BEG2;
	output S1BEG3;
	output S2BEG0;
	output S2BEG1;
	output S2BEG2;
	output S2BEG3;
	output S2BEG4;
	output S2BEG5;
	output S2BEG6;
	output S2BEG7;
	output S2BEGb0;
	output S2BEGb1;
	output S2BEGb2;
	output S2BEGb3;
	output S2BEGb4;
	output S2BEGb5;
	output S2BEGb6;
	output S2BEGb7;
	output S4BEG0;
	output S4BEG1;
	output S4BEG2;
	output S4BEG3;
	output W1BEG0;
	output W1BEG1;
	output W1BEG2;
	output W1BEG3;
	output W2BEG0;
	output W2BEG1;
	output W2BEG2;
	output W2BEG3;
	output W2BEG4;
	output W2BEG5;
	output W2BEG6;
	output W2BEG7;
	output W2BEGb0;
	output W2BEGb1;
	output W2BEGb2;
	output W2BEGb3;
	output W2BEGb4;
	output W2BEGb5;
	output W2BEGb6;
	output W2BEGb7;
	output WW4BEG0;
	output WW4BEG1;
	output WW4BEG2;
	output WW4BEG3;
	output WW4BEG4;
	output WW4BEG5;
	output WW4BEG6;
	output WW4BEG7;
	output WW4BEG8;
	output WW4BEG9;
	output WW4BEG10;
	output WW4BEG11;
	output WW4BEG12;
	output WW4BEG13;
	output WW4BEG14;
	output WW4BEG15;
	output W6BEG0;
	output W6BEG1;
	output W6BEG2;
	output W6BEG3;
	output W6BEG4;
	output W6BEG5;
	output W6BEG6;
	output W6BEG7;
	output W6BEG8;
	output W6BEG9;
	output W6BEG10;
	output W6BEG11;
	output FAB2RAM_D0_I0;
	output FAB2RAM_D0_I1;
	output FAB2RAM_D0_I2;
	output FAB2RAM_D0_I3;
	output FAB2RAM_D1_I0;
	output FAB2RAM_D1_I1;
	output FAB2RAM_D1_I2;
	output FAB2RAM_D1_I3;
	output FAB2RAM_D2_I0;
	output FAB2RAM_D2_I1;
	output FAB2RAM_D2_I2;
	output FAB2RAM_D2_I3;
	output FAB2RAM_D3_I0;
	output FAB2RAM_D3_I1;
	output FAB2RAM_D3_I2;
	output FAB2RAM_D3_I3;
	output FAB2RAM_A0_I0;
	output FAB2RAM_A0_I1;
	output FAB2RAM_A0_I2;
	output FAB2RAM_A0_I3;
	output FAB2RAM_A1_I0;
	output FAB2RAM_A1_I1;
	output FAB2RAM_A1_I2;
	output FAB2RAM_A1_I3;
	output FAB2RAM_C_I0;
	output FAB2RAM_C_I1;
	output FAB2RAM_C_I2;
	output FAB2RAM_C_I3;
	output J_NS4_BEG0;
	output J_NS4_BEG1;
	output J_NS4_BEG2;
	output J_NS4_BEG3;
	output J_NS4_BEG4;
	output J_NS4_BEG5;
	output J_NS4_BEG6;
	output J_NS4_BEG7;
	output J_NS4_BEG8;
	output J_NS4_BEG9;
	output J_NS4_BEG10;
	output J_NS4_BEG11;
	output J_NS4_BEG12;
	output J_NS4_BEG13;
	output J_NS4_BEG14;
	output J_NS4_BEG15;
	output J_NS2_BEG0;
	output J_NS2_BEG1;
	output J_NS2_BEG2;
	output J_NS2_BEG3;
	output J_NS2_BEG4;
	output J_NS2_BEG5;
	output J_NS2_BEG6;
	output J_NS2_BEG7;
	output J_NS1_BEG0;
	output J_NS1_BEG1;
	output J_NS1_BEG2;
	output J_NS1_BEG3;
	//global
	input [NoConfigBits-1:0] ConfigBits;
	input [NoConfigBits-1:0] ConfigBits_N;

	parameter GND0 = 1'b0;
	parameter GND = 1'b0;
	parameter VCC0 = 1'b1;
	parameter VCC = 1'b1;
	parameter VDD0 = 1'b1;
	parameter VDD = 1'b1;
	
	wire [4-1:0] N1BEG0_input;
	wire [4-1:0] N1BEG1_input;
	wire [4-1:0] N1BEG2_input;
	wire [4-1:0] N1BEG3_input;
	wire [4-1:0] N2BEG0_input;
	wire [4-1:0] N2BEG1_input;
	wire [4-1:0] N2BEG2_input;
	wire [4-1:0] N2BEG3_input;
	wire [4-1:0] N2BEG4_input;
	wire [4-1:0] N2BEG5_input;
	wire [4-1:0] N2BEG6_input;
	wire [4-1:0] N2BEG7_input;
	wire [1-1:0] N2BEGb0_input;
	wire [1-1:0] N2BEGb1_input;
	wire [1-1:0] N2BEGb2_input;
	wire [1-1:0] N2BEGb3_input;
	wire [1-1:0] N2BEGb4_input;
	wire [1-1:0] N2BEGb5_input;
	wire [1-1:0] N2BEGb6_input;
	wire [1-1:0] N2BEGb7_input;
	wire [8-1:0] N4BEG0_input;
	wire [8-1:0] N4BEG1_input;
	wire [8-1:0] N4BEG2_input;
	wire [8-1:0] N4BEG3_input;
	wire [4-1:0] S1BEG0_input;
	wire [4-1:0] S1BEG1_input;
	wire [4-1:0] S1BEG2_input;
	wire [4-1:0] S1BEG3_input;
	wire [4-1:0] S2BEG0_input;
	wire [4-1:0] S2BEG1_input;
	wire [4-1:0] S2BEG2_input;
	wire [4-1:0] S2BEG3_input;
	wire [4-1:0] S2BEG4_input;
	wire [4-1:0] S2BEG5_input;
	wire [4-1:0] S2BEG6_input;
	wire [4-1:0] S2BEG7_input;
	wire [1-1:0] S2BEGb0_input;
	wire [1-1:0] S2BEGb1_input;
	wire [1-1:0] S2BEGb2_input;
	wire [1-1:0] S2BEGb3_input;
	wire [1-1:0] S2BEGb4_input;
	wire [1-1:0] S2BEGb5_input;
	wire [1-1:0] S2BEGb6_input;
	wire [1-1:0] S2BEGb7_input;
	wire [8-1:0] S4BEG0_input;
	wire [8-1:0] S4BEG1_input;
	wire [8-1:0] S4BEG2_input;
	wire [8-1:0] S4BEG3_input;
	wire [4-1:0] W1BEG0_input;
	wire [4-1:0] W1BEG1_input;
	wire [4-1:0] W1BEG2_input;
	wire [4-1:0] W1BEG3_input;
	wire [4-1:0] W2BEG0_input;
	wire [4-1:0] W2BEG1_input;
	wire [4-1:0] W2BEG2_input;
	wire [4-1:0] W2BEG3_input;
	wire [4-1:0] W2BEG4_input;
	wire [4-1:0] W2BEG5_input;
	wire [4-1:0] W2BEG6_input;
	wire [4-1:0] W2BEG7_input;
	wire [4-1:0] W2BEGb0_input;
	wire [4-1:0] W2BEGb1_input;
	wire [4-1:0] W2BEGb2_input;
	wire [4-1:0] W2BEGb3_input;
	wire [4-1:0] W2BEGb4_input;
	wire [4-1:0] W2BEGb5_input;
	wire [4-1:0] W2BEGb6_input;
	wire [4-1:0] W2BEGb7_input;
	wire [4-1:0] WW4BEG0_input;
	wire [4-1:0] WW4BEG1_input;
	wire [4-1:0] WW4BEG2_input;
	wire [4-1:0] WW4BEG3_input;
	wire [4-1:0] WW4BEG4_input;
	wire [4-1:0] WW4BEG5_input;
	wire [4-1:0] WW4BEG6_input;
	wire [4-1:0] WW4BEG7_input;
	wire [4-1:0] WW4BEG8_input;
	wire [4-1:0] WW4BEG9_input;
	wire [4-1:0] WW4BEG10_input;
	wire [4-1:0] WW4BEG11_input;
	wire [4-1:0] WW4BEG12_input;
	wire [4-1:0] WW4BEG13_input;
	wire [4-1:0] WW4BEG14_input;
	wire [4-1:0] WW4BEG15_input;
	wire [4-1:0] W6BEG0_input;
	wire [4-1:0] W6BEG1_input;
	wire [4-1:0] W6BEG2_input;
	wire [4-1:0] W6BEG3_input;
	wire [4-1:0] W6BEG4_input;
	wire [4-1:0] W6BEG5_input;
	wire [4-1:0] W6BEG6_input;
	wire [4-1:0] W6BEG7_input;
	wire [4-1:0] W6BEG8_input;
	wire [4-1:0] W6BEG9_input;
	wire [4-1:0] W6BEG10_input;
	wire [4-1:0] W6BEG11_input;
	wire [4-1:0] FAB2RAM_D0_I0_input;
	wire [4-1:0] FAB2RAM_D0_I1_input;
	wire [4-1:0] FAB2RAM_D0_I2_input;
	wire [4-1:0] FAB2RAM_D0_I3_input;
	wire [4-1:0] FAB2RAM_D1_I0_input;
	wire [4-1:0] FAB2RAM_D1_I1_input;
	wire [4-1:0] FAB2RAM_D1_I2_input;
	wire [4-1:0] FAB2RAM_D1_I3_input;
	wire [4-1:0] FAB2RAM_D2_I0_input;
	wire [4-1:0] FAB2RAM_D2_I1_input;
	wire [4-1:0] FAB2RAM_D2_I2_input;
	wire [4-1:0] FAB2RAM_D2_I3_input;
	wire [4-1:0] FAB2RAM_D3_I0_input;
	wire [4-1:0] FAB2RAM_D3_I1_input;
	wire [4-1:0] FAB2RAM_D3_I2_input;
	wire [4-1:0] FAB2RAM_D3_I3_input;
	wire [4-1:0] FAB2RAM_A0_I0_input;
	wire [4-1:0] FAB2RAM_A0_I1_input;
	wire [4-1:0] FAB2RAM_A0_I2_input;
	wire [4-1:0] FAB2RAM_A0_I3_input;
	wire [4-1:0] FAB2RAM_A1_I0_input;
	wire [4-1:0] FAB2RAM_A1_I1_input;
	wire [4-1:0] FAB2RAM_A1_I2_input;
	wire [4-1:0] FAB2RAM_A1_I3_input;
	wire [4-1:0] FAB2RAM_C_I0_input;
	wire [4-1:0] FAB2RAM_C_I1_input;
	wire [4-1:0] FAB2RAM_C_I2_input;
	wire [4-1:0] FAB2RAM_C_I3_input;
	wire [4-1:0] J_NS4_BEG0_input;
	wire [4-1:0] J_NS4_BEG1_input;
	wire [4-1:0] J_NS4_BEG2_input;
	wire [4-1:0] J_NS4_BEG3_input;
	wire [4-1:0] J_NS4_BEG4_input;
	wire [4-1:0] J_NS4_BEG5_input;
	wire [4-1:0] J_NS4_BEG6_input;
	wire [4-1:0] J_NS4_BEG7_input;
	wire [4-1:0] J_NS4_BEG8_input;
	wire [4-1:0] J_NS4_BEG9_input;
	wire [4-1:0] J_NS4_BEG10_input;
	wire [4-1:0] J_NS4_BEG11_input;
	wire [4-1:0] J_NS4_BEG12_input;
	wire [4-1:0] J_NS4_BEG13_input;
	wire [4-1:0] J_NS4_BEG14_input;
	wire [4-1:0] J_NS4_BEG15_input;
	wire [4-1:0] J_NS2_BEG0_input;
	wire [4-1:0] J_NS2_BEG1_input;
	wire [4-1:0] J_NS2_BEG2_input;
	wire [4-1:0] J_NS2_BEG3_input;
	wire [4-1:0] J_NS2_BEG4_input;
	wire [4-1:0] J_NS2_BEG5_input;
	wire [4-1:0] J_NS2_BEG6_input;
	wire [4-1:0] J_NS2_BEG7_input;
	wire [4-1:0] J_NS1_BEG0_input;
	wire [4-1:0] J_NS1_BEG1_input;
	wire [4-1:0] J_NS1_BEG2_input;
	wire [4-1:0] J_NS1_BEG3_input;

	wire [2-1:0] DEBUG_select_N1BEG0;
	wire [2-1:0] DEBUG_select_N1BEG1;
	wire [2-1:0] DEBUG_select_N1BEG2;
	wire [2-1:0] DEBUG_select_N1BEG3;
	wire [2-1:0] DEBUG_select_N2BEG0;
	wire [2-1:0] DEBUG_select_N2BEG1;
	wire [2-1:0] DEBUG_select_N2BEG2;
	wire [2-1:0] DEBUG_select_N2BEG3;
	wire [2-1:0] DEBUG_select_N2BEG4;
	wire [2-1:0] DEBUG_select_N2BEG5;
	wire [2-1:0] DEBUG_select_N2BEG6;
	wire [2-1:0] DEBUG_select_N2BEG7;
	wire [3-1:0] DEBUG_select_N4BEG0;
	wire [3-1:0] DEBUG_select_N4BEG1;
	wire [3-1:0] DEBUG_select_N4BEG2;
	wire [3-1:0] DEBUG_select_N4BEG3;
	wire [2-1:0] DEBUG_select_S1BEG0;
	wire [2-1:0] DEBUG_select_S1BEG1;
	wire [2-1:0] DEBUG_select_S1BEG2;
	wire [2-1:0] DEBUG_select_S1BEG3;
	wire [2-1:0] DEBUG_select_S2BEG0;
	wire [2-1:0] DEBUG_select_S2BEG1;
	wire [2-1:0] DEBUG_select_S2BEG2;
	wire [2-1:0] DEBUG_select_S2BEG3;
	wire [2-1:0] DEBUG_select_S2BEG4;
	wire [2-1:0] DEBUG_select_S2BEG5;
	wire [2-1:0] DEBUG_select_S2BEG6;
	wire [2-1:0] DEBUG_select_S2BEG7;
	wire [3-1:0] DEBUG_select_S4BEG0;
	wire [3-1:0] DEBUG_select_S4BEG1;
	wire [3-1:0] DEBUG_select_S4BEG2;
	wire [3-1:0] DEBUG_select_S4BEG3;
	wire [2-1:0] DEBUG_select_W1BEG0;
	wire [2-1:0] DEBUG_select_W1BEG1;
	wire [2-1:0] DEBUG_select_W1BEG2;
	wire [2-1:0] DEBUG_select_W1BEG3;
	wire [2-1:0] DEBUG_select_W2BEG0;
	wire [2-1:0] DEBUG_select_W2BEG1;
	wire [2-1:0] DEBUG_select_W2BEG2;
	wire [2-1:0] DEBUG_select_W2BEG3;
	wire [2-1:0] DEBUG_select_W2BEG4;
	wire [2-1:0] DEBUG_select_W2BEG5;
	wire [2-1:0] DEBUG_select_W2BEG6;
	wire [2-1:0] DEBUG_select_W2BEG7;
	wire [2-1:0] DEBUG_select_W2BEGb0;
	wire [2-1:0] DEBUG_select_W2BEGb1;
	wire [2-1:0] DEBUG_select_W2BEGb2;
	wire [2-1:0] DEBUG_select_W2BEGb3;
	wire [2-1:0] DEBUG_select_W2BEGb4;
	wire [2-1:0] DEBUG_select_W2BEGb5;
	wire [2-1:0] DEBUG_select_W2BEGb6;
	wire [2-1:0] DEBUG_select_W2BEGb7;
	wire [2-1:0] DEBUG_select_WW4BEG0;
	wire [2-1:0] DEBUG_select_WW4BEG1;
	wire [2-1:0] DEBUG_select_WW4BEG2;
	wire [2-1:0] DEBUG_select_WW4BEG3;
	wire [2-1:0] DEBUG_select_WW4BEG4;
	wire [2-1:0] DEBUG_select_WW4BEG5;
	wire [2-1:0] DEBUG_select_WW4BEG6;
	wire [2-1:0] DEBUG_select_WW4BEG7;
	wire [2-1:0] DEBUG_select_WW4BEG8;
	wire [2-1:0] DEBUG_select_WW4BEG9;
	wire [2-1:0] DEBUG_select_WW4BEG10;
	wire [2-1:0] DEBUG_select_WW4BEG11;
	wire [2-1:0] DEBUG_select_WW4BEG12;
	wire [2-1:0] DEBUG_select_WW4BEG13;
	wire [2-1:0] DEBUG_select_WW4BEG14;
	wire [2-1:0] DEBUG_select_WW4BEG15;
	wire [2-1:0] DEBUG_select_W6BEG0;
	wire [2-1:0] DEBUG_select_W6BEG1;
	wire [2-1:0] DEBUG_select_W6BEG2;
	wire [2-1:0] DEBUG_select_W6BEG3;
	wire [2-1:0] DEBUG_select_W6BEG4;
	wire [2-1:0] DEBUG_select_W6BEG5;
	wire [2-1:0] DEBUG_select_W6BEG6;
	wire [2-1:0] DEBUG_select_W6BEG7;
	wire [2-1:0] DEBUG_select_W6BEG8;
	wire [2-1:0] DEBUG_select_W6BEG9;
	wire [2-1:0] DEBUG_select_W6BEG10;
	wire [2-1:0] DEBUG_select_W6BEG11;
	wire [2-1:0] DEBUG_select_FAB2RAM_D0_I0;
	wire [2-1:0] DEBUG_select_FAB2RAM_D0_I1;
	wire [2-1:0] DEBUG_select_FAB2RAM_D0_I2;
	wire [2-1:0] DEBUG_select_FAB2RAM_D0_I3;
	wire [2-1:0] DEBUG_select_FAB2RAM_D1_I0;
	wire [2-1:0] DEBUG_select_FAB2RAM_D1_I1;
	wire [2-1:0] DEBUG_select_FAB2RAM_D1_I2;
	wire [2-1:0] DEBUG_select_FAB2RAM_D1_I3;
	wire [2-1:0] DEBUG_select_FAB2RAM_D2_I0;
	wire [2-1:0] DEBUG_select_FAB2RAM_D2_I1;
	wire [2-1:0] DEBUG_select_FAB2RAM_D2_I2;
	wire [2-1:0] DEBUG_select_FAB2RAM_D2_I3;
	wire [2-1:0] DEBUG_select_FAB2RAM_D3_I0;
	wire [2-1:0] DEBUG_select_FAB2RAM_D3_I1;
	wire [2-1:0] DEBUG_select_FAB2RAM_D3_I2;
	wire [2-1:0] DEBUG_select_FAB2RAM_D3_I3;
	wire [2-1:0] DEBUG_select_FAB2RAM_A0_I0;
	wire [2-1:0] DEBUG_select_FAB2RAM_A0_I1;
	wire [2-1:0] DEBUG_select_FAB2RAM_A0_I2;
	wire [2-1:0] DEBUG_select_FAB2RAM_A0_I3;
	wire [2-1:0] DEBUG_select_FAB2RAM_A1_I0;
	wire [2-1:0] DEBUG_select_FAB2RAM_A1_I1;
	wire [2-1:0] DEBUG_select_FAB2RAM_A1_I2;
	wire [2-1:0] DEBUG_select_FAB2RAM_A1_I3;
	wire [2-1:0] DEBUG_select_FAB2RAM_C_I0;
	wire [2-1:0] DEBUG_select_FAB2RAM_C_I1;
	wire [2-1:0] DEBUG_select_FAB2RAM_C_I2;
	wire [2-1:0] DEBUG_select_FAB2RAM_C_I3;
	wire [2-1:0] DEBUG_select_J_NS4_BEG0;
	wire [2-1:0] DEBUG_select_J_NS4_BEG1;
	wire [2-1:0] DEBUG_select_J_NS4_BEG2;
	wire [2-1:0] DEBUG_select_J_NS4_BEG3;
	wire [2-1:0] DEBUG_select_J_NS4_BEG4;
	wire [2-1:0] DEBUG_select_J_NS4_BEG5;
	wire [2-1:0] DEBUG_select_J_NS4_BEG6;
	wire [2-1:0] DEBUG_select_J_NS4_BEG7;
	wire [2-1:0] DEBUG_select_J_NS4_BEG8;
	wire [2-1:0] DEBUG_select_J_NS4_BEG9;
	wire [2-1:0] DEBUG_select_J_NS4_BEG10;
	wire [2-1:0] DEBUG_select_J_NS4_BEG11;
	wire [2-1:0] DEBUG_select_J_NS4_BEG12;
	wire [2-1:0] DEBUG_select_J_NS4_BEG13;
	wire [2-1:0] DEBUG_select_J_NS4_BEG14;
	wire [2-1:0] DEBUG_select_J_NS4_BEG15;
	wire [2-1:0] DEBUG_select_J_NS2_BEG0;
	wire [2-1:0] DEBUG_select_J_NS2_BEG1;
	wire [2-1:0] DEBUG_select_J_NS2_BEG2;
	wire [2-1:0] DEBUG_select_J_NS2_BEG3;
	wire [2-1:0] DEBUG_select_J_NS2_BEG4;
	wire [2-1:0] DEBUG_select_J_NS2_BEG5;
	wire [2-1:0] DEBUG_select_J_NS2_BEG6;
	wire [2-1:0] DEBUG_select_J_NS2_BEG7;
	wire [2-1:0] DEBUG_select_J_NS1_BEG0;
	wire [2-1:0] DEBUG_select_J_NS1_BEG1;
	wire [2-1:0] DEBUG_select_J_NS1_BEG2;
	wire [2-1:0] DEBUG_select_J_NS1_BEG3;

// The configuration bits (if any) are just a long shift register

// This shift register is padded to an even number of flops/latches
// switch matrix multiplexer  N1BEG0 		MUX-4
	assign N1BEG0_input = {J_NS1_END0,J_NS4_END12,E6END4,E1END0};
	assign N1BEG0 = N1BEG0_input[ConfigBits[1:0]];
 
// switch matrix multiplexer  N1BEG1 		MUX-4
	assign N1BEG1_input = {J_NS1_END1,J_NS4_END13,E6END5,E1END1};
	assign N1BEG1 = N1BEG1_input[ConfigBits[3:2]];
 
// switch matrix multiplexer  N1BEG2 		MUX-4
	assign N1BEG2_input = {J_NS1_END2,J_NS4_END14,E6END6,E1END2};
	assign N1BEG2 = N1BEG2_input[ConfigBits[5:4]];
 
// switch matrix multiplexer  N1BEG3 		MUX-4
	assign N1BEG3_input = {J_NS1_END3,J_NS4_END15,E6END7,E1END3};
	assign N1BEG3 = N1BEG3_input[ConfigBits[7:6]];
 
// switch matrix multiplexer  N2BEG0 		MUX-4
	assign N2BEG0_input = {J_NS2_END0,E6END7,E2END7,E2MID7};
	assign N2BEG0 = N2BEG0_input[ConfigBits[9:8]];
 
// switch matrix multiplexer  N2BEG1 		MUX-4
	assign N2BEG1_input = {J_NS2_END1,E6END6,E2END6,E2MID6};
	assign N2BEG1 = N2BEG1_input[ConfigBits[11:10]];
 
// switch matrix multiplexer  N2BEG2 		MUX-4
	assign N2BEG2_input = {J_NS2_END2,E6END5,E2END5,E2MID5};
	assign N2BEG2 = N2BEG2_input[ConfigBits[13:12]];
 
// switch matrix multiplexer  N2BEG3 		MUX-4
	assign N2BEG3_input = {J_NS2_END3,E6END4,E2END4,E2MID4};
	assign N2BEG3 = N2BEG3_input[ConfigBits[15:14]];
 
// switch matrix multiplexer  N2BEG4 		MUX-4
	assign N2BEG4_input = {J_NS2_END4,E6END3,E2END3,E2MID3};
	assign N2BEG4 = N2BEG4_input[ConfigBits[17:16]];
 
// switch matrix multiplexer  N2BEG5 		MUX-4
	assign N2BEG5_input = {J_NS2_END5,E6END2,E2END2,E2MID2};
	assign N2BEG5 = N2BEG5_input[ConfigBits[19:18]];
 
// switch matrix multiplexer  N2BEG6 		MUX-4
	assign N2BEG6_input = {J_NS2_END6,E6END1,E2END1,E2MID1};
	assign N2BEG6 = N2BEG6_input[ConfigBits[21:20]];
 
// switch matrix multiplexer  N2BEG7 		MUX-4
	assign N2BEG7_input = {J_NS2_END7,E6END0,E2END0,E2MID0};
	assign N2BEG7 = N2BEG7_input[ConfigBits[23:22]];
 
// switch matrix multiplexer  N2BEGb0 		MUX-1
	assign N2BEGb0 = N2MID0;
// switch matrix multiplexer  N2BEGb1 		MUX-1
	assign N2BEGb1 = N2MID1;
// switch matrix multiplexer  N2BEGb2 		MUX-1
	assign N2BEGb2 = N2MID2;
// switch matrix multiplexer  N2BEGb3 		MUX-1
	assign N2BEGb3 = N2MID3;
// switch matrix multiplexer  N2BEGb4 		MUX-1
	assign N2BEGb4 = N2MID4;
// switch matrix multiplexer  N2BEGb5 		MUX-1
	assign N2BEGb5 = N2MID5;
// switch matrix multiplexer  N2BEGb6 		MUX-1
	assign N2BEGb6 = N2MID6;
// switch matrix multiplexer  N2BEGb7 		MUX-1
	assign N2BEGb7 = N2MID7;
// switch matrix multiplexer  N4BEG0 		MUX-8
	assign N4BEG0_input = {J_NS2_END0,J_NS4_END12,J_NS4_END8,J_NS4_END4,J_NS4_END0,E6END8,EE4END0,E1END0};
	assign N4BEG0 = N4BEG0_input[ConfigBits[26:24]];
 
// switch matrix multiplexer  N4BEG1 		MUX-8
	assign N4BEG1_input = {J_NS2_END1,J_NS4_END13,J_NS4_END9,J_NS4_END5,J_NS4_END1,E6END9,EE4END1,E1END1};
	assign N4BEG1 = N4BEG1_input[ConfigBits[29:27]];
 
// switch matrix multiplexer  N4BEG2 		MUX-8
	assign N4BEG2_input = {J_NS2_END2,J_NS4_END14,J_NS4_END10,J_NS4_END6,J_NS4_END2,E6END10,EE4END2,E1END2};
	assign N4BEG2 = N4BEG2_input[ConfigBits[32:30]];
 
// switch matrix multiplexer  N4BEG3 		MUX-8
	assign N4BEG3_input = {J_NS2_END3,J_NS4_END15,J_NS4_END11,J_NS4_END7,J_NS4_END3,E6END11,EE4END3,E1END3};
	assign N4BEG3 = N4BEG3_input[ConfigBits[35:33]];
 
// switch matrix multiplexer  S1BEG0 		MUX-4
	assign S1BEG0_input = {J_NS1_END0,J_NS4_END12,E6END8,E1END0};
	assign S1BEG0 = S1BEG0_input[ConfigBits[37:36]];
 
// switch matrix multiplexer  S1BEG1 		MUX-4
	assign S1BEG1_input = {J_NS1_END1,J_NS4_END13,E6END9,E1END1};
	assign S1BEG1 = S1BEG1_input[ConfigBits[39:38]];
 
// switch matrix multiplexer  S1BEG2 		MUX-4
	assign S1BEG2_input = {J_NS1_END2,J_NS4_END14,E6END10,E1END2};
	assign S1BEG2 = S1BEG2_input[ConfigBits[41:40]];
 
// switch matrix multiplexer  S1BEG3 		MUX-4
	assign S1BEG3_input = {J_NS1_END3,J_NS4_END15,E6END11,E1END3};
	assign S1BEG3 = S1BEG3_input[ConfigBits[43:42]];
 
// switch matrix multiplexer  S2BEG0 		MUX-4
	assign S2BEG0_input = {J_NS2_END0,E6END8,E2END7,E2MID7};
	assign S2BEG0 = S2BEG0_input[ConfigBits[45:44]];
 
// switch matrix multiplexer  S2BEG1 		MUX-4
	assign S2BEG1_input = {J_NS2_END1,E6END9,E2END6,E2MID6};
	assign S2BEG1 = S2BEG1_input[ConfigBits[47:46]];
 
// switch matrix multiplexer  S2BEG2 		MUX-4
	assign S2BEG2_input = {J_NS2_END2,E6END10,E2END5,E2MID5};
	assign S2BEG2 = S2BEG2_input[ConfigBits[49:48]];
 
// switch matrix multiplexer  S2BEG3 		MUX-4
	assign S2BEG3_input = {J_NS2_END3,E6END11,E2END4,E2MID4};
	assign S2BEG3 = S2BEG3_input[ConfigBits[51:50]];
 
// switch matrix multiplexer  S2BEG4 		MUX-4
	assign S2BEG4_input = {J_NS2_END4,E2END3,E2MID3,E1END0};
	assign S2BEG4 = S2BEG4_input[ConfigBits[53:52]];
 
// switch matrix multiplexer  S2BEG5 		MUX-4
	assign S2BEG5_input = {J_NS2_END5,E2END2,E2MID2,E1END1};
	assign S2BEG5 = S2BEG5_input[ConfigBits[55:54]];
 
// switch matrix multiplexer  S2BEG6 		MUX-4
	assign S2BEG6_input = {J_NS2_END6,E2END1,E2MID1,E1END2};
	assign S2BEG6 = S2BEG6_input[ConfigBits[57:56]];
 
// switch matrix multiplexer  S2BEG7 		MUX-4
	assign S2BEG7_input = {J_NS2_END7,E2END0,E2MID0,E1END3};
	assign S2BEG7 = S2BEG7_input[ConfigBits[59:58]];
 
// switch matrix multiplexer  S2BEGb0 		MUX-1
	assign S2BEGb0 = S2MID0;
// switch matrix multiplexer  S2BEGb1 		MUX-1
	assign S2BEGb1 = S2MID1;
// switch matrix multiplexer  S2BEGb2 		MUX-1
	assign S2BEGb2 = S2MID2;
// switch matrix multiplexer  S2BEGb3 		MUX-1
	assign S2BEGb3 = S2MID3;
// switch matrix multiplexer  S2BEGb4 		MUX-1
	assign S2BEGb4 = S2MID4;
// switch matrix multiplexer  S2BEGb5 		MUX-1
	assign S2BEGb5 = S2MID5;
// switch matrix multiplexer  S2BEGb6 		MUX-1
	assign S2BEGb6 = S2MID6;
// switch matrix multiplexer  S2BEGb7 		MUX-1
	assign S2BEGb7 = S2MID7;
// switch matrix multiplexer  S4BEG0 		MUX-8
	assign S4BEG0_input = {J_NS2_END4,J_NS4_END12,J_NS4_END8,J_NS4_END4,J_NS4_END0,E6END4,EE4END12,E1END0};
	assign S4BEG0 = S4BEG0_input[ConfigBits[62:60]];
 
// switch matrix multiplexer  S4BEG1 		MUX-8
	assign S4BEG1_input = {J_NS2_END5,J_NS4_END13,J_NS4_END9,J_NS4_END5,J_NS4_END1,E6END5,EE4END13,E1END1};
	assign S4BEG1 = S4BEG1_input[ConfigBits[65:63]];
 
// switch matrix multiplexer  S4BEG2 		MUX-8
	assign S4BEG2_input = {J_NS2_END6,J_NS4_END14,J_NS4_END10,J_NS4_END6,J_NS4_END2,E6END6,EE4END14,E1END2};
	assign S4BEG2 = S4BEG2_input[ConfigBits[68:66]];
 
// switch matrix multiplexer  S4BEG3 		MUX-8
	assign S4BEG3_input = {J_NS2_END7,J_NS4_END15,J_NS4_END11,J_NS4_END7,J_NS4_END3,E6END7,EE4END15,E1END3};
	assign S4BEG3 = S4BEG3_input[ConfigBits[71:69]];
 
// switch matrix multiplexer  W1BEG0 		MUX-4
	assign W1BEG0_input = {RAM2FAB_D1_O3,RAM2FAB_D0_O2,S1END0,N1END0};
	assign W1BEG0 = W1BEG0_input[ConfigBits[73:72]];
 
// switch matrix multiplexer  W1BEG1 		MUX-4
	assign W1BEG1_input = {RAM2FAB_D1_O2,RAM2FAB_D0_O3,S1END1,N1END1};
	assign W1BEG1 = W1BEG1_input[ConfigBits[75:74]];
 
// switch matrix multiplexer  W1BEG2 		MUX-4
	assign W1BEG2_input = {RAM2FAB_D1_O1,RAM2FAB_D0_O0,S1END2,N1END2};
	assign W1BEG2 = W1BEG2_input[ConfigBits[77:76]];
 
// switch matrix multiplexer  W1BEG3 		MUX-4
	assign W1BEG3_input = {RAM2FAB_D1_O0,RAM2FAB_D0_O1,S1END3,N1END3};
	assign W1BEG3 = W1BEG3_input[ConfigBits[79:78]];
 
// switch matrix multiplexer  W2BEG0 		MUX-4
	assign W2BEG0_input = {J_NS2_END7,J_NS2_END0,RAM2FAB_D2_O0,RAM2FAB_D0_O0};
	assign W2BEG0 = W2BEG0_input[ConfigBits[81:80]];
 
// switch matrix multiplexer  W2BEG1 		MUX-4
	assign W2BEG1_input = {J_NS2_END6,J_NS2_END1,RAM2FAB_D2_O1,RAM2FAB_D0_O1};
	assign W2BEG1 = W2BEG1_input[ConfigBits[83:82]];
 
// switch matrix multiplexer  W2BEG2 		MUX-4
	assign W2BEG2_input = {J_NS2_END5,J_NS2_END2,RAM2FAB_D2_O2,RAM2FAB_D0_O2};
	assign W2BEG2 = W2BEG2_input[ConfigBits[85:84]];
 
// switch matrix multiplexer  W2BEG3 		MUX-4
	assign W2BEG3_input = {J_NS2_END4,J_NS2_END3,RAM2FAB_D2_O3,RAM2FAB_D0_O3};
	assign W2BEG3 = W2BEG3_input[ConfigBits[87:86]];
 
// switch matrix multiplexer  W2BEG4 		MUX-4
	assign W2BEG4_input = {J_NS2_END4,J_NS2_END3,RAM2FAB_D3_O0,RAM2FAB_D1_O0};
	assign W2BEG4 = W2BEG4_input[ConfigBits[89:88]];
 
// switch matrix multiplexer  W2BEG5 		MUX-4
	assign W2BEG5_input = {J_NS2_END5,J_NS2_END2,RAM2FAB_D3_O1,RAM2FAB_D1_O1};
	assign W2BEG5 = W2BEG5_input[ConfigBits[91:90]];
 
// switch matrix multiplexer  W2BEG6 		MUX-4
	assign W2BEG6_input = {J_NS2_END6,J_NS2_END1,RAM2FAB_D3_O2,RAM2FAB_D1_O2};
	assign W2BEG6 = W2BEG6_input[ConfigBits[93:92]];
 
// switch matrix multiplexer  W2BEG7 		MUX-4
	assign W2BEG7_input = {J_NS2_END7,J_NS2_END0,RAM2FAB_D3_O3,RAM2FAB_D1_O3};
	assign W2BEG7 = W2BEG7_input[ConfigBits[95:94]];
 
// switch matrix multiplexer  W2BEGb0 		MUX-4
	assign W2BEGb0_input = {J_NS2_END7,J_NS2_END0,RAM2FAB_D2_O0,RAM2FAB_D0_O0};
	assign W2BEGb0 = W2BEGb0_input[ConfigBits[97:96]];
 
// switch matrix multiplexer  W2BEGb1 		MUX-4
	assign W2BEGb1_input = {J_NS2_END6,J_NS2_END1,RAM2FAB_D2_O1,RAM2FAB_D0_O1};
	assign W2BEGb1 = W2BEGb1_input[ConfigBits[99:98]];
 
// switch matrix multiplexer  W2BEGb2 		MUX-4
	assign W2BEGb2_input = {J_NS2_END5,J_NS2_END2,RAM2FAB_D2_O2,RAM2FAB_D0_O2};
	assign W2BEGb2 = W2BEGb2_input[ConfigBits[101:100]];
 
// switch matrix multiplexer  W2BEGb3 		MUX-4
	assign W2BEGb3_input = {J_NS2_END4,J_NS2_END3,RAM2FAB_D2_O3,RAM2FAB_D0_O3};
	assign W2BEGb3 = W2BEGb3_input[ConfigBits[103:102]];
 
// switch matrix multiplexer  W2BEGb4 		MUX-4
	assign W2BEGb4_input = {J_NS2_END4,J_NS2_END3,RAM2FAB_D3_O0,RAM2FAB_D1_O0};
	assign W2BEGb4 = W2BEGb4_input[ConfigBits[105:104]];
 
// switch matrix multiplexer  W2BEGb5 		MUX-4
	assign W2BEGb5_input = {J_NS2_END5,J_NS2_END2,RAM2FAB_D3_O1,RAM2FAB_D1_O1};
	assign W2BEGb5 = W2BEGb5_input[ConfigBits[107:106]];
 
// switch matrix multiplexer  W2BEGb6 		MUX-4
	assign W2BEGb6_input = {J_NS2_END6,J_NS2_END1,RAM2FAB_D3_O2,RAM2FAB_D1_O2};
	assign W2BEGb6 = W2BEGb6_input[ConfigBits[109:108]];
 
// switch matrix multiplexer  W2BEGb7 		MUX-4
	assign W2BEGb7_input = {J_NS2_END7,J_NS2_END0,RAM2FAB_D3_O3,RAM2FAB_D1_O3};
	assign W2BEGb7 = W2BEGb7_input[ConfigBits[111:110]];
 
// switch matrix multiplexer  WW4BEG0 		MUX-4
	assign WW4BEG0_input = {J_NS2_END7,J_NS4_END15,RAM2FAB_D3_O0,RAM2FAB_D0_O0};
	assign WW4BEG0 = WW4BEG0_input[ConfigBits[113:112]];
 
// switch matrix multiplexer  WW4BEG1 		MUX-4
	assign WW4BEG1_input = {J_NS2_END6,J_NS4_END14,RAM2FAB_D3_O1,RAM2FAB_D0_O1};
	assign WW4BEG1 = WW4BEG1_input[ConfigBits[115:114]];
 
// switch matrix multiplexer  WW4BEG2 		MUX-4
	assign WW4BEG2_input = {J_NS2_END5,J_NS4_END13,RAM2FAB_D3_O2,RAM2FAB_D0_O2};
	assign WW4BEG2 = WW4BEG2_input[ConfigBits[117:116]];
 
// switch matrix multiplexer  WW4BEG3 		MUX-4
	assign WW4BEG3_input = {J_NS2_END4,J_NS4_END12,RAM2FAB_D3_O3,RAM2FAB_D0_O3};
	assign WW4BEG3 = WW4BEG3_input[ConfigBits[119:118]];
 
// switch matrix multiplexer  WW4BEG4 		MUX-4
	assign WW4BEG4_input = {J_NS2_END3,J_NS4_END11,RAM2FAB_D2_O0,RAM2FAB_D1_O0};
	assign WW4BEG4 = WW4BEG4_input[ConfigBits[121:120]];
 
// switch matrix multiplexer  WW4BEG5 		MUX-4
	assign WW4BEG5_input = {J_NS2_END2,J_NS4_END10,RAM2FAB_D2_O1,RAM2FAB_D1_O1};
	assign WW4BEG5 = WW4BEG5_input[ConfigBits[123:122]];
 
// switch matrix multiplexer  WW4BEG6 		MUX-4
	assign WW4BEG6_input = {J_NS2_END1,J_NS4_END9,RAM2FAB_D2_O2,RAM2FAB_D1_O2};
	assign WW4BEG6 = WW4BEG6_input[ConfigBits[125:124]];
 
// switch matrix multiplexer  WW4BEG7 		MUX-4
	assign WW4BEG7_input = {J_NS2_END0,J_NS4_END8,RAM2FAB_D2_O3,RAM2FAB_D1_O3};
	assign WW4BEG7 = WW4BEG7_input[ConfigBits[127:126]];
 
// switch matrix multiplexer  WW4BEG8 		MUX-4
	assign WW4BEG8_input = {J_NS2_END7,J_NS4_END7,RAM2FAB_D2_O0,RAM2FAB_D1_O0};
	assign WW4BEG8 = WW4BEG8_input[ConfigBits[129:128]];
 
// switch matrix multiplexer  WW4BEG9 		MUX-4
	assign WW4BEG9_input = {J_NS2_END6,J_NS4_END6,RAM2FAB_D2_O1,RAM2FAB_D1_O1};
	assign WW4BEG9 = WW4BEG9_input[ConfigBits[131:130]];
 
// switch matrix multiplexer  WW4BEG10 		MUX-4
	assign WW4BEG10_input = {J_NS2_END5,J_NS4_END5,RAM2FAB_D2_O2,RAM2FAB_D1_O2};
	assign WW4BEG10 = WW4BEG10_input[ConfigBits[133:132]];
 
// switch matrix multiplexer  WW4BEG11 		MUX-4
	assign WW4BEG11_input = {J_NS2_END4,J_NS4_END4,RAM2FAB_D2_O3,RAM2FAB_D1_O3};
	assign WW4BEG11 = WW4BEG11_input[ConfigBits[135:134]];
 
// switch matrix multiplexer  WW4BEG12 		MUX-4
	assign WW4BEG12_input = {J_NS2_END3,J_NS4_END3,RAM2FAB_D3_O0,RAM2FAB_D0_O0};
	assign WW4BEG12 = WW4BEG12_input[ConfigBits[137:136]];
 
// switch matrix multiplexer  WW4BEG13 		MUX-4
	assign WW4BEG13_input = {J_NS2_END2,J_NS4_END2,RAM2FAB_D3_O1,RAM2FAB_D0_O1};
	assign WW4BEG13 = WW4BEG13_input[ConfigBits[139:138]];
 
// switch matrix multiplexer  WW4BEG14 		MUX-4
	assign WW4BEG14_input = {J_NS2_END1,J_NS4_END1,RAM2FAB_D3_O2,RAM2FAB_D0_O2};
	assign WW4BEG14 = WW4BEG14_input[ConfigBits[141:140]];
 
// switch matrix multiplexer  WW4BEG15 		MUX-4
	assign WW4BEG15_input = {J_NS2_END0,J_NS4_END0,RAM2FAB_D3_O3,RAM2FAB_D0_O3};
	assign WW4BEG15 = WW4BEG15_input[ConfigBits[143:142]];
 
// switch matrix multiplexer  W6BEG0 		MUX-4
	assign W6BEG0_input = {J_NS4_END15,J_NS4_END11,S4END0,N4END0};
	assign W6BEG0 = W6BEG0_input[ConfigBits[145:144]];
 
// switch matrix multiplexer  W6BEG1 		MUX-4
	assign W6BEG1_input = {J_NS4_END14,J_NS4_END10,S4END1,N4END1};
	assign W6BEG1 = W6BEG1_input[ConfigBits[147:146]];
 
// switch matrix multiplexer  W6BEG2 		MUX-4
	assign W6BEG2_input = {J_NS4_END13,J_NS4_END9,S4END2,N4END2};
	assign W6BEG2 = W6BEG2_input[ConfigBits[149:148]];
 
// switch matrix multiplexer  W6BEG3 		MUX-4
	assign W6BEG3_input = {J_NS4_END12,J_NS4_END8,S4END3,N4END3};
	assign W6BEG3 = W6BEG3_input[ConfigBits[151:150]];
 
// switch matrix multiplexer  W6BEG4 		MUX-4
	assign W6BEG4_input = {J_NS2_END0,J_NS4_END11,J_NS4_END7,RAM2FAB_D1_O0};
	assign W6BEG4 = W6BEG4_input[ConfigBits[153:152]];
 
// switch matrix multiplexer  W6BEG5 		MUX-4
	assign W6BEG5_input = {J_NS2_END1,J_NS4_END10,J_NS4_END6,RAM2FAB_D1_O1};
	assign W6BEG5 = W6BEG5_input[ConfigBits[155:154]];
 
// switch matrix multiplexer  W6BEG6 		MUX-4
	assign W6BEG6_input = {J_NS2_END2,J_NS4_END9,J_NS4_END5,RAM2FAB_D1_O2};
	assign W6BEG6 = W6BEG6_input[ConfigBits[157:156]];
 
// switch matrix multiplexer  W6BEG7 		MUX-4
	assign W6BEG7_input = {J_NS2_END3,J_NS4_END8,J_NS4_END4,RAM2FAB_D1_O3};
	assign W6BEG7 = W6BEG7_input[ConfigBits[159:158]];
 
// switch matrix multiplexer  W6BEG8 		MUX-4
	assign W6BEG8_input = {J_NS2_END4,J_NS4_END7,J_NS4_END3,RAM2FAB_D0_O0};
	assign W6BEG8 = W6BEG8_input[ConfigBits[161:160]];
 
// switch matrix multiplexer  W6BEG9 		MUX-4
	assign W6BEG9_input = {J_NS2_END5,J_NS4_END6,J_NS4_END2,RAM2FAB_D0_O1};
	assign W6BEG9 = W6BEG9_input[ConfigBits[163:162]];
 
// switch matrix multiplexer  W6BEG10 		MUX-4
	assign W6BEG10_input = {J_NS2_END6,J_NS4_END5,J_NS4_END1,RAM2FAB_D0_O2};
	assign W6BEG10 = W6BEG10_input[ConfigBits[165:164]];
 
// switch matrix multiplexer  W6BEG11 		MUX-4
	assign W6BEG11_input = {J_NS2_END7,J_NS4_END4,J_NS4_END0,RAM2FAB_D0_O3};
	assign W6BEG11 = W6BEG11_input[ConfigBits[167:166]];
 
// switch matrix multiplexer  FAB2RAM_D0_I0 		MUX-4
	assign FAB2RAM_D0_I0_input = {J_NS4_END0,E6END0,EE4END8,EE4END0};
	assign FAB2RAM_D0_I0 = FAB2RAM_D0_I0_input[ConfigBits[169:168]];
 
// switch matrix multiplexer  FAB2RAM_D0_I1 		MUX-4
	assign FAB2RAM_D0_I1_input = {J_NS4_END1,E6END1,EE4END9,EE4END1};
	assign FAB2RAM_D0_I1 = FAB2RAM_D0_I1_input[ConfigBits[171:170]];
 
// switch matrix multiplexer  FAB2RAM_D0_I2 		MUX-4
	assign FAB2RAM_D0_I2_input = {J_NS4_END2,E6END2,EE4END10,EE4END2};
	assign FAB2RAM_D0_I2 = FAB2RAM_D0_I2_input[ConfigBits[173:172]];
 
// switch matrix multiplexer  FAB2RAM_D0_I3 		MUX-4
	assign FAB2RAM_D0_I3_input = {J_NS4_END3,E6END3,EE4END11,EE4END3};
	assign FAB2RAM_D0_I3 = FAB2RAM_D0_I3_input[ConfigBits[175:174]];
 
// switch matrix multiplexer  FAB2RAM_D1_I0 		MUX-4
	assign FAB2RAM_D1_I0_input = {J_NS4_END4,E6END4,EE4END12,EE4END4};
	assign FAB2RAM_D1_I0 = FAB2RAM_D1_I0_input[ConfigBits[177:176]];
 
// switch matrix multiplexer  FAB2RAM_D1_I1 		MUX-4
	assign FAB2RAM_D1_I1_input = {J_NS4_END5,E6END5,EE4END13,EE4END5};
	assign FAB2RAM_D1_I1 = FAB2RAM_D1_I1_input[ConfigBits[179:178]];
 
// switch matrix multiplexer  FAB2RAM_D1_I2 		MUX-4
	assign FAB2RAM_D1_I2_input = {J_NS4_END6,E6END6,EE4END14,EE4END6};
	assign FAB2RAM_D1_I2 = FAB2RAM_D1_I2_input[ConfigBits[181:180]];
 
// switch matrix multiplexer  FAB2RAM_D1_I3 		MUX-4
	assign FAB2RAM_D1_I3_input = {J_NS4_END7,E6END7,EE4END15,EE4END7};
	assign FAB2RAM_D1_I3 = FAB2RAM_D1_I3_input[ConfigBits[183:182]];
 
// switch matrix multiplexer  FAB2RAM_D2_I0 		MUX-4
	assign FAB2RAM_D2_I0_input = {J_NS4_END8,E6END8,EE4END8,EE4END0};
	assign FAB2RAM_D2_I0 = FAB2RAM_D2_I0_input[ConfigBits[185:184]];
 
// switch matrix multiplexer  FAB2RAM_D2_I1 		MUX-4
	assign FAB2RAM_D2_I1_input = {J_NS4_END9,E6END9,EE4END9,EE4END1};
	assign FAB2RAM_D2_I1 = FAB2RAM_D2_I1_input[ConfigBits[187:186]];
 
// switch matrix multiplexer  FAB2RAM_D2_I2 		MUX-4
	assign FAB2RAM_D2_I2_input = {J_NS4_END10,E6END10,EE4END10,EE4END2};
	assign FAB2RAM_D2_I2 = FAB2RAM_D2_I2_input[ConfigBits[189:188]];
 
// switch matrix multiplexer  FAB2RAM_D2_I3 		MUX-4
	assign FAB2RAM_D2_I3_input = {J_NS4_END11,E6END11,EE4END11,EE4END3};
	assign FAB2RAM_D2_I3 = FAB2RAM_D2_I3_input[ConfigBits[191:190]];
 
// switch matrix multiplexer  FAB2RAM_D3_I0 		MUX-4
	assign FAB2RAM_D3_I0_input = {J_NS4_END12,EE4END12,EE4END4,E1END0};
	assign FAB2RAM_D3_I0 = FAB2RAM_D3_I0_input[ConfigBits[193:192]];
 
// switch matrix multiplexer  FAB2RAM_D3_I1 		MUX-4
	assign FAB2RAM_D3_I1_input = {J_NS4_END13,EE4END13,EE4END5,E1END1};
	assign FAB2RAM_D3_I1 = FAB2RAM_D3_I1_input[ConfigBits[195:194]];
 
// switch matrix multiplexer  FAB2RAM_D3_I2 		MUX-4
	assign FAB2RAM_D3_I2_input = {J_NS4_END14,EE4END14,EE4END6,E1END2};
	assign FAB2RAM_D3_I2 = FAB2RAM_D3_I2_input[ConfigBits[197:196]];
 
// switch matrix multiplexer  FAB2RAM_D3_I3 		MUX-4
	assign FAB2RAM_D3_I3_input = {J_NS4_END15,EE4END15,EE4END7,E1END3};
	assign FAB2RAM_D3_I3 = FAB2RAM_D3_I3_input[ConfigBits[199:198]];
 
// switch matrix multiplexer  FAB2RAM_A0_I0 		MUX-4
	assign FAB2RAM_A0_I0_input = {GND0,J_NS2_END0,E2END0,E2MID0};
	assign FAB2RAM_A0_I0 = FAB2RAM_A0_I0_input[ConfigBits[201:200]];
 
// switch matrix multiplexer  FAB2RAM_A0_I1 		MUX-4
	assign FAB2RAM_A0_I1_input = {GND0,J_NS2_END1,E2END1,E2MID1};
	assign FAB2RAM_A0_I1 = FAB2RAM_A0_I1_input[ConfigBits[203:202]];
 
// switch matrix multiplexer  FAB2RAM_A0_I2 		MUX-4
	assign FAB2RAM_A0_I2_input = {GND0,J_NS2_END2,E2END2,E2MID2};
	assign FAB2RAM_A0_I2 = FAB2RAM_A0_I2_input[ConfigBits[205:204]];
 
// switch matrix multiplexer  FAB2RAM_A0_I3 		MUX-4
	assign FAB2RAM_A0_I3_input = {GND0,J_NS2_END3,E2END3,E2MID3};
	assign FAB2RAM_A0_I3 = FAB2RAM_A0_I3_input[ConfigBits[207:206]];
 
// switch matrix multiplexer  FAB2RAM_A1_I0 		MUX-4
	assign FAB2RAM_A1_I0_input = {GND0,J_NS2_END4,E2END4,E2MID4};
	assign FAB2RAM_A1_I0 = FAB2RAM_A1_I0_input[ConfigBits[209:208]];
 
// switch matrix multiplexer  FAB2RAM_A1_I1 		MUX-4
	assign FAB2RAM_A1_I1_input = {GND0,J_NS2_END5,E2END5,E2MID5};
	assign FAB2RAM_A1_I1 = FAB2RAM_A1_I1_input[ConfigBits[211:210]];
 
// switch matrix multiplexer  FAB2RAM_A1_I2 		MUX-4
	assign FAB2RAM_A1_I2_input = {GND0,J_NS2_END6,E2END6,E2MID6};
	assign FAB2RAM_A1_I2 = FAB2RAM_A1_I2_input[ConfigBits[213:212]];
 
// switch matrix multiplexer  FAB2RAM_A1_I3 		MUX-4
	assign FAB2RAM_A1_I3_input = {GND0,J_NS2_END7,E2END7,E2MID7};
	assign FAB2RAM_A1_I3 = FAB2RAM_A1_I3_input[ConfigBits[215:214]];
 
// switch matrix multiplexer  FAB2RAM_C_I0 		MUX-4
	assign FAB2RAM_C_I0_input = {GND0,J_NS1_END0,E6END0,E1END0};
	assign FAB2RAM_C_I0 = FAB2RAM_C_I0_input[ConfigBits[217:216]];
 
// switch matrix multiplexer  FAB2RAM_C_I1 		MUX-4
	assign FAB2RAM_C_I1_input = {GND0,J_NS1_END1,E6END1,E1END1};
	assign FAB2RAM_C_I1 = FAB2RAM_C_I1_input[ConfigBits[219:218]];
 
// switch matrix multiplexer  FAB2RAM_C_I2 		MUX-4
	assign FAB2RAM_C_I2_input = {GND0,J_NS1_END2,E6END2,E1END2};
	assign FAB2RAM_C_I2 = FAB2RAM_C_I2_input[ConfigBits[221:220]];
 
// switch matrix multiplexer  FAB2RAM_C_I3 		MUX-4
	assign FAB2RAM_C_I3_input = {GND0,J_NS1_END3,E6END3,E1END3};
	assign FAB2RAM_C_I3 = FAB2RAM_C_I3_input[ConfigBits[223:222]];
 
// switch matrix multiplexer  J_NS4_BEG0 		MUX-4
	assign J_NS4_BEG0_input = {S4END0,S1END0,N4END0,N1END0};
	assign J_NS4_BEG0 = J_NS4_BEG0_input[ConfigBits[225:224]];
 
// switch matrix multiplexer  J_NS4_BEG1 		MUX-4
	assign J_NS4_BEG1_input = {S4END1,S1END1,N4END1,N1END1};
	assign J_NS4_BEG1 = J_NS4_BEG1_input[ConfigBits[227:226]];
 
// switch matrix multiplexer  J_NS4_BEG2 		MUX-4
	assign J_NS4_BEG2_input = {S4END2,S1END2,N4END2,N1END2};
	assign J_NS4_BEG2 = J_NS4_BEG2_input[ConfigBits[229:228]];
 
// switch matrix multiplexer  J_NS4_BEG3 		MUX-4
	assign J_NS4_BEG3_input = {S4END3,S1END3,N4END3,N1END3};
	assign J_NS4_BEG3 = J_NS4_BEG3_input[ConfigBits[231:230]];
 
// switch matrix multiplexer  J_NS4_BEG4 		MUX-4
	assign J_NS4_BEG4_input = {S4END0,S1END0,N4END0,N1END0};
	assign J_NS4_BEG4 = J_NS4_BEG4_input[ConfigBits[233:232]];
 
// switch matrix multiplexer  J_NS4_BEG5 		MUX-4
	assign J_NS4_BEG5_input = {S4END1,S1END1,N4END1,N1END1};
	assign J_NS4_BEG5 = J_NS4_BEG5_input[ConfigBits[235:234]];
 
// switch matrix multiplexer  J_NS4_BEG6 		MUX-4
	assign J_NS4_BEG6_input = {S4END2,S1END2,N4END2,N1END2};
	assign J_NS4_BEG6 = J_NS4_BEG6_input[ConfigBits[237:236]];
 
// switch matrix multiplexer  J_NS4_BEG7 		MUX-4
	assign J_NS4_BEG7_input = {S4END3,S1END3,N4END3,N1END3};
	assign J_NS4_BEG7 = J_NS4_BEG7_input[ConfigBits[239:238]];
 
// switch matrix multiplexer  J_NS4_BEG8 		MUX-4
	assign J_NS4_BEG8_input = {S4END0,S1END0,N4END0,N1END0};
	assign J_NS4_BEG8 = J_NS4_BEG8_input[ConfigBits[241:240]];
 
// switch matrix multiplexer  J_NS4_BEG9 		MUX-4
	assign J_NS4_BEG9_input = {S4END1,S1END1,N4END1,N1END1};
	assign J_NS4_BEG9 = J_NS4_BEG9_input[ConfigBits[243:242]];
 
// switch matrix multiplexer  J_NS4_BEG10 		MUX-4
	assign J_NS4_BEG10_input = {S4END2,S1END2,N4END2,N1END2};
	assign J_NS4_BEG10 = J_NS4_BEG10_input[ConfigBits[245:244]];
 
// switch matrix multiplexer  J_NS4_BEG11 		MUX-4
	assign J_NS4_BEG11_input = {S4END3,S1END3,N4END3,N1END3};
	assign J_NS4_BEG11 = J_NS4_BEG11_input[ConfigBits[247:246]];
 
// switch matrix multiplexer  J_NS4_BEG12 		MUX-4
	assign J_NS4_BEG12_input = {S4END0,S1END0,N4END0,N1END0};
	assign J_NS4_BEG12 = J_NS4_BEG12_input[ConfigBits[249:248]];
 
// switch matrix multiplexer  J_NS4_BEG13 		MUX-4
	assign J_NS4_BEG13_input = {S4END1,S1END1,N4END1,N1END1};
	assign J_NS4_BEG13 = J_NS4_BEG13_input[ConfigBits[251:250]];
 
// switch matrix multiplexer  J_NS4_BEG14 		MUX-4
	assign J_NS4_BEG14_input = {S4END2,S1END2,N4END2,N1END2};
	assign J_NS4_BEG14 = J_NS4_BEG14_input[ConfigBits[253:252]];
 
// switch matrix multiplexer  J_NS4_BEG15 		MUX-4
	assign J_NS4_BEG15_input = {S4END3,S1END3,N4END3,N1END3};
	assign J_NS4_BEG15 = J_NS4_BEG15_input[ConfigBits[255:254]];
 
// switch matrix multiplexer  J_NS2_BEG0 		MUX-4
	assign J_NS2_BEG0_input = {S2END0,S2MID0,N2END0,N2MID0};
	assign J_NS2_BEG0 = J_NS2_BEG0_input[ConfigBits[257:256]];
 
// switch matrix multiplexer  J_NS2_BEG1 		MUX-4
	assign J_NS2_BEG1_input = {S2END1,S2MID1,N2END1,N2MID1};
	assign J_NS2_BEG1 = J_NS2_BEG1_input[ConfigBits[259:258]];
 
// switch matrix multiplexer  J_NS2_BEG2 		MUX-4
	assign J_NS2_BEG2_input = {S2END2,S2MID2,N2END2,N2MID2};
	assign J_NS2_BEG2 = J_NS2_BEG2_input[ConfigBits[261:260]];
 
// switch matrix multiplexer  J_NS2_BEG3 		MUX-4
	assign J_NS2_BEG3_input = {S2END3,S2MID3,N2END3,N2MID3};
	assign J_NS2_BEG3 = J_NS2_BEG3_input[ConfigBits[263:262]];
 
// switch matrix multiplexer  J_NS2_BEG4 		MUX-4
	assign J_NS2_BEG4_input = {S2END4,S2MID4,N2END4,N2MID4};
	assign J_NS2_BEG4 = J_NS2_BEG4_input[ConfigBits[265:264]];
 
// switch matrix multiplexer  J_NS2_BEG5 		MUX-4
	assign J_NS2_BEG5_input = {S2END5,S2MID5,N2END5,N2MID5};
	assign J_NS2_BEG5 = J_NS2_BEG5_input[ConfigBits[267:266]];
 
// switch matrix multiplexer  J_NS2_BEG6 		MUX-4
	assign J_NS2_BEG6_input = {S2END6,S2MID6,N2END6,N2MID6};
	assign J_NS2_BEG6 = J_NS2_BEG6_input[ConfigBits[269:268]];
 
// switch matrix multiplexer  J_NS2_BEG7 		MUX-4
	assign J_NS2_BEG7_input = {S2END7,S2MID7,N2END7,N2MID7};
	assign J_NS2_BEG7 = J_NS2_BEG7_input[ConfigBits[271:270]];
 
// switch matrix multiplexer  J_NS1_BEG0 		MUX-4
	assign J_NS1_BEG0_input = {GND0,S1END0,E6END0,N1END0};
	assign J_NS1_BEG0 = J_NS1_BEG0_input[ConfigBits[273:272]];
 
// switch matrix multiplexer  J_NS1_BEG1 		MUX-4
	assign J_NS1_BEG1_input = {GND0,S1END1,E6END1,N1END1};
	assign J_NS1_BEG1 = J_NS1_BEG1_input[ConfigBits[275:274]];
 
// switch matrix multiplexer  J_NS1_BEG2 		MUX-4
	assign J_NS1_BEG2_input = {GND0,S1END2,E6END2,N1END2};
	assign J_NS1_BEG2 = J_NS1_BEG2_input[ConfigBits[277:276]];
 
// switch matrix multiplexer  J_NS1_BEG3 		MUX-4
	assign J_NS1_BEG3_input = {GND0,S1END3,E6END3,N1END3};
	assign J_NS1_BEG3 = J_NS1_BEG3_input[ConfigBits[279:278]];
 
	assign DEBUG_select_N1BEG0 = ConfigBits[1:0];
	assign DEBUG_select_N1BEG1 = ConfigBits[3:2];
	assign DEBUG_select_N1BEG2 = ConfigBits[5:4];
	assign DEBUG_select_N1BEG3 = ConfigBits[7:6];
	assign DEBUG_select_N2BEG0 = ConfigBits[9:8];
	assign DEBUG_select_N2BEG1 = ConfigBits[11:10];
	assign DEBUG_select_N2BEG2 = ConfigBits[13:12];
	assign DEBUG_select_N2BEG3 = ConfigBits[15:14];
	assign DEBUG_select_N2BEG4 = ConfigBits[17:16];
	assign DEBUG_select_N2BEG5 = ConfigBits[19:18];
	assign DEBUG_select_N2BEG6 = ConfigBits[21:20];
	assign DEBUG_select_N2BEG7 = ConfigBits[23:22];
	assign DEBUG_select_N4BEG0 = ConfigBits[26:24];
	assign DEBUG_select_N4BEG1 = ConfigBits[29:27];
	assign DEBUG_select_N4BEG2 = ConfigBits[32:30];
	assign DEBUG_select_N4BEG3 = ConfigBits[35:33];
	assign DEBUG_select_S1BEG0 = ConfigBits[37:36];
	assign DEBUG_select_S1BEG1 = ConfigBits[39:38];
	assign DEBUG_select_S1BEG2 = ConfigBits[41:40];
	assign DEBUG_select_S1BEG3 = ConfigBits[43:42];
	assign DEBUG_select_S2BEG0 = ConfigBits[45:44];
	assign DEBUG_select_S2BEG1 = ConfigBits[47:46];
	assign DEBUG_select_S2BEG2 = ConfigBits[49:48];
	assign DEBUG_select_S2BEG3 = ConfigBits[51:50];
	assign DEBUG_select_S2BEG4 = ConfigBits[53:52];
	assign DEBUG_select_S2BEG5 = ConfigBits[55:54];
	assign DEBUG_select_S2BEG6 = ConfigBits[57:56];
	assign DEBUG_select_S2BEG7 = ConfigBits[59:58];
	assign DEBUG_select_S4BEG0 = ConfigBits[62:60];
	assign DEBUG_select_S4BEG1 = ConfigBits[65:63];
	assign DEBUG_select_S4BEG2 = ConfigBits[68:66];
	assign DEBUG_select_S4BEG3 = ConfigBits[71:69];
	assign DEBUG_select_W1BEG0 = ConfigBits[73:72];
	assign DEBUG_select_W1BEG1 = ConfigBits[75:74];
	assign DEBUG_select_W1BEG2 = ConfigBits[77:76];
	assign DEBUG_select_W1BEG3 = ConfigBits[79:78];
	assign DEBUG_select_W2BEG0 = ConfigBits[81:80];
	assign DEBUG_select_W2BEG1 = ConfigBits[83:82];
	assign DEBUG_select_W2BEG2 = ConfigBits[85:84];
	assign DEBUG_select_W2BEG3 = ConfigBits[87:86];
	assign DEBUG_select_W2BEG4 = ConfigBits[89:88];
	assign DEBUG_select_W2BEG5 = ConfigBits[91:90];
	assign DEBUG_select_W2BEG6 = ConfigBits[93:92];
	assign DEBUG_select_W2BEG7 = ConfigBits[95:94];
	assign DEBUG_select_W2BEGb0 = ConfigBits[97:96];
	assign DEBUG_select_W2BEGb1 = ConfigBits[99:98];
	assign DEBUG_select_W2BEGb2 = ConfigBits[101:100];
	assign DEBUG_select_W2BEGb3 = ConfigBits[103:102];
	assign DEBUG_select_W2BEGb4 = ConfigBits[105:104];
	assign DEBUG_select_W2BEGb5 = ConfigBits[107:106];
	assign DEBUG_select_W2BEGb6 = ConfigBits[109:108];
	assign DEBUG_select_W2BEGb7 = ConfigBits[111:110];
	assign DEBUG_select_WW4BEG0 = ConfigBits[113:112];
	assign DEBUG_select_WW4BEG1 = ConfigBits[115:114];
	assign DEBUG_select_WW4BEG2 = ConfigBits[117:116];
	assign DEBUG_select_WW4BEG3 = ConfigBits[119:118];
	assign DEBUG_select_WW4BEG4 = ConfigBits[121:120];
	assign DEBUG_select_WW4BEG5 = ConfigBits[123:122];
	assign DEBUG_select_WW4BEG6 = ConfigBits[125:124];
	assign DEBUG_select_WW4BEG7 = ConfigBits[127:126];
	assign DEBUG_select_WW4BEG8 = ConfigBits[129:128];
	assign DEBUG_select_WW4BEG9 = ConfigBits[131:130];
	assign DEBUG_select_WW4BEG10 = ConfigBits[133:132];
	assign DEBUG_select_WW4BEG11 = ConfigBits[135:134];
	assign DEBUG_select_WW4BEG12 = ConfigBits[137:136];
	assign DEBUG_select_WW4BEG13 = ConfigBits[139:138];
	assign DEBUG_select_WW4BEG14 = ConfigBits[141:140];
	assign DEBUG_select_WW4BEG15 = ConfigBits[143:142];
	assign DEBUG_select_W6BEG0 = ConfigBits[145:144];
	assign DEBUG_select_W6BEG1 = ConfigBits[147:146];
	assign DEBUG_select_W6BEG2 = ConfigBits[149:148];
	assign DEBUG_select_W6BEG3 = ConfigBits[151:150];
	assign DEBUG_select_W6BEG4 = ConfigBits[153:152];
	assign DEBUG_select_W6BEG5 = ConfigBits[155:154];
	assign DEBUG_select_W6BEG6 = ConfigBits[157:156];
	assign DEBUG_select_W6BEG7 = ConfigBits[159:158];
	assign DEBUG_select_W6BEG8 = ConfigBits[161:160];
	assign DEBUG_select_W6BEG9 = ConfigBits[163:162];
	assign DEBUG_select_W6BEG10 = ConfigBits[165:164];
	assign DEBUG_select_W6BEG11 = ConfigBits[167:166];
	assign DEBUG_select_FAB2RAM_D0_I0 = ConfigBits[169:168];
	assign DEBUG_select_FAB2RAM_D0_I1 = ConfigBits[171:170];
	assign DEBUG_select_FAB2RAM_D0_I2 = ConfigBits[173:172];
	assign DEBUG_select_FAB2RAM_D0_I3 = ConfigBits[175:174];
	assign DEBUG_select_FAB2RAM_D1_I0 = ConfigBits[177:176];
	assign DEBUG_select_FAB2RAM_D1_I1 = ConfigBits[179:178];
	assign DEBUG_select_FAB2RAM_D1_I2 = ConfigBits[181:180];
	assign DEBUG_select_FAB2RAM_D1_I3 = ConfigBits[183:182];
	assign DEBUG_select_FAB2RAM_D2_I0 = ConfigBits[185:184];
	assign DEBUG_select_FAB2RAM_D2_I1 = ConfigBits[187:186];
	assign DEBUG_select_FAB2RAM_D2_I2 = ConfigBits[189:188];
	assign DEBUG_select_FAB2RAM_D2_I3 = ConfigBits[191:190];
	assign DEBUG_select_FAB2RAM_D3_I0 = ConfigBits[193:192];
	assign DEBUG_select_FAB2RAM_D3_I1 = ConfigBits[195:194];
	assign DEBUG_select_FAB2RAM_D3_I2 = ConfigBits[197:196];
	assign DEBUG_select_FAB2RAM_D3_I3 = ConfigBits[199:198];
	assign DEBUG_select_FAB2RAM_A0_I0 = ConfigBits[201:200];
	assign DEBUG_select_FAB2RAM_A0_I1 = ConfigBits[203:202];
	assign DEBUG_select_FAB2RAM_A0_I2 = ConfigBits[205:204];
	assign DEBUG_select_FAB2RAM_A0_I3 = ConfigBits[207:206];
	assign DEBUG_select_FAB2RAM_A1_I0 = ConfigBits[209:208];
	assign DEBUG_select_FAB2RAM_A1_I1 = ConfigBits[211:210];
	assign DEBUG_select_FAB2RAM_A1_I2 = ConfigBits[213:212];
	assign DEBUG_select_FAB2RAM_A1_I3 = ConfigBits[215:214];
	assign DEBUG_select_FAB2RAM_C_I0 = ConfigBits[217:216];
	assign DEBUG_select_FAB2RAM_C_I1 = ConfigBits[219:218];
	assign DEBUG_select_FAB2RAM_C_I2 = ConfigBits[221:220];
	assign DEBUG_select_FAB2RAM_C_I3 = ConfigBits[223:222];
	assign DEBUG_select_J_NS4_BEG0 = ConfigBits[225:224];
	assign DEBUG_select_J_NS4_BEG1 = ConfigBits[227:226];
	assign DEBUG_select_J_NS4_BEG2 = ConfigBits[229:228];
	assign DEBUG_select_J_NS4_BEG3 = ConfigBits[231:230];
	assign DEBUG_select_J_NS4_BEG4 = ConfigBits[233:232];
	assign DEBUG_select_J_NS4_BEG5 = ConfigBits[235:234];
	assign DEBUG_select_J_NS4_BEG6 = ConfigBits[237:236];
	assign DEBUG_select_J_NS4_BEG7 = ConfigBits[239:238];
	assign DEBUG_select_J_NS4_BEG8 = ConfigBits[241:240];
	assign DEBUG_select_J_NS4_BEG9 = ConfigBits[243:242];
	assign DEBUG_select_J_NS4_BEG10 = ConfigBits[245:244];
	assign DEBUG_select_J_NS4_BEG11 = ConfigBits[247:246];
	assign DEBUG_select_J_NS4_BEG12 = ConfigBits[249:248];
	assign DEBUG_select_J_NS4_BEG13 = ConfigBits[251:250];
	assign DEBUG_select_J_NS4_BEG14 = ConfigBits[253:252];
	assign DEBUG_select_J_NS4_BEG15 = ConfigBits[255:254];
	assign DEBUG_select_J_NS2_BEG0 = ConfigBits[257:256];
	assign DEBUG_select_J_NS2_BEG1 = ConfigBits[259:258];
	assign DEBUG_select_J_NS2_BEG2 = ConfigBits[261:260];
	assign DEBUG_select_J_NS2_BEG3 = ConfigBits[263:262];
	assign DEBUG_select_J_NS2_BEG4 = ConfigBits[265:264];
	assign DEBUG_select_J_NS2_BEG5 = ConfigBits[267:266];
	assign DEBUG_select_J_NS2_BEG6 = ConfigBits[269:268];
	assign DEBUG_select_J_NS2_BEG7 = ConfigBits[271:270];
	assign DEBUG_select_J_NS1_BEG0 = ConfigBits[273:272];
	assign DEBUG_select_J_NS1_BEG1 = ConfigBits[275:274];
	assign DEBUG_select_J_NS1_BEG2 = ConfigBits[277:276];
	assign DEBUG_select_J_NS1_BEG3 = ConfigBits[279:278];

endmodule
